module Module58();
    Module77 inst_Module77();
endmodule
