module rootModule_sub0_0_sub1_2();
    rootModule_sub0_0_sub1_2_sub2_0 inst_0();
    rootModule_sub0_0_sub1_2_sub2_1 inst_1();
endmodule
