module Module81();
    Module97 inst_Module97();
    Module87 inst_Module87();
    Module91 inst_Module91();
    Module82 inst_Module82();
endmodule
