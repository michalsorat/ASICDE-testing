module rootModule_2_2_1_0_1();
endmodule
