module Module38();
    Module83 inst_Module83();
    Module71 inst_Module71();
endmodule
