module Module3();
    Module56 inst_Module56();
    Module94 inst_Module94();
    Module15 inst_Module15();
endmodule
