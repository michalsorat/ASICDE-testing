module rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_2_se7_0_se8_3();
    rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_2_se7_0_se8_3_se9_0 inst_0();
    rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_2_se7_0_se8_3_se9_1 inst_1();
    rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_2_se7_0_se8_3_se9_2 inst_2();
    rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_2_se7_0_se8_3_se9_3 inst_3();
    rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_2_se7_0_se8_3_se9_4 inst_4();
endmodule
