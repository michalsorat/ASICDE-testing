module Module26();
    Module58 inst_Module58();
    Module73 inst_Module73();
    Module59 inst_Module59();
endmodule
