module rootModule_sub0_0_sub1_1();
    rootModule_sub0_0_sub1_1_sub2_0 inst_0();
    rootModule_sub0_0_sub1_1_sub2_1 inst_1();
    rootModule_sub0_0_sub1_1_sub2_2 inst_2();
endmodule
