module rootModule_sb0_0_sb1_1_sb2_2_sb3_1_sb4_1();
endmodule
