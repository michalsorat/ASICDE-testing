module rootModule_sub0_0_sub1_0_sub2_1_sub3_1_sub4_2();
endmodule
