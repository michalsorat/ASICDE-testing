module Module56();
    Module70 inst_Module70();
    Module89 inst_Module89();
    Module90 inst_Module90();
    Module74 inst_Module74();
    Module71 inst_Module71();
endmodule
