module rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_1_sw7_0_sw8_4_sw9_4();
endmodule
