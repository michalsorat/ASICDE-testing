module rootModule_2_1_0_0_0();
endmodule
