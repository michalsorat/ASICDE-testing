module rootModule_1_1_0_0_0();
endmodule
