module rootModule_sb0_1_sb1_1_sb2_2();
    rootModule_sb0_1_sb1_1_sb2_2_sb3_0 inst_0();
    rootModule_sb0_1_sb1_1_sb2_2_sb3_1 inst_1();
    rootModule_sb0_1_sb1_1_sb2_2_sb3_2 inst_2();
endmodule
