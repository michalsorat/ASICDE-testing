module rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0();
    rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0 inst_0();
endmodule
