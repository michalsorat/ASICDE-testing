module rootModule_sub_0_1_sub_1_0_sub_2_2_sub_3_1();
    rootModule_sub_0_1_sub_1_0_sub_2_2_sub_3_1_sub_4_0 inst_0();
    rootModule_sub_0_1_sub_1_0_sub_2_2_sub_3_1_sub_4_1 inst_1();
    rootModule_sub_0_1_sub_1_0_sub_2_2_sub_3_1_sub_4_2 inst_2();
endmodule
