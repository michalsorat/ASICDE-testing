module rootModule_sb0_0_sb1_2_sb2_1_sb3_2_sb4_2();
endmodule
