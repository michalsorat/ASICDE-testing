module rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_0_sg8_2();
    rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_0_sg8_2_sg9_0 inst_0();
    rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_0_sg8_2_sg9_1 inst_1();
    rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_0_sg8_2_sg9_2 inst_2();
    rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_0_sg8_2_sg9_3 inst_3();
    rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_0_sg8_2_sg9_4 inst_4();
endmodule
