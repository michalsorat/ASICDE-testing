module Module93();
    Module98 inst_Module98();
    Module97 inst_Module97();
endmodule
