module rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_0_sc7_1_sc8_2_sc9_2();
endmodule
