module Module51();
    Module88 inst_Module88();
    Module89 inst_Module89();
    Module65 inst_Module65();
    Module72 inst_Module72();
    Module76 inst_Module76();
endmodule
