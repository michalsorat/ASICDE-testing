module Module16();
    Module34 inst_Module34();
    Module78 inst_Module78();
    Module17 inst_Module17();
endmodule
