module Module57();
    Module93 inst_Module93();
    Module97 inst_Module97();
    Module61 inst_Module61();
endmodule
