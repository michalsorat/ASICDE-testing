module rootModule_1_0_0_0_0();
endmodule
