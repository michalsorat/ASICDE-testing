module rootModule_sb0_1_sb1_2_sb2_1_sb3_1_sb4_1();
endmodule
