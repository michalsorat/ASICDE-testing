module rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0();
    rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0 inst_0();
endmodule
