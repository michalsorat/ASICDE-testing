module rootModule_sub0_0();
    rootModule_sub0_0_sub1_0 inst_0();
endmodule
