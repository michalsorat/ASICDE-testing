module Module1();
    Module35 inst_Module35();
    Module81 inst_Module81();
    Module42 inst_Module42();
    Module73 inst_Module73();
endmodule
