module Module30();
    Module35 inst_Module35();
    Module76 inst_Module76();
    Module56 inst_Module56();
    Module62 inst_Module62();
endmodule
