module rootModule_sb0_0_sb1_2();
    rootModule_sb0_0_sb1_2_sb2_0 inst_0();
    rootModule_sb0_0_sb1_2_sb2_1 inst_1();
    rootModule_sb0_0_sb1_2_sb2_2 inst_2();
endmodule
