module rootModule_sg0_0_sg1_0();
    rootModule_sg0_0_sg1_0_sg2_0 inst_0();
endmodule
