module Module32();
    Module53 inst_Module53();
    Module91 inst_Module91();
    Module76 inst_Module76();
    Module44 inst_Module44();
    Module55 inst_Module55();
endmodule
