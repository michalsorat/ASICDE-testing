module Module24();
    Module45 inst_Module45();
    Module70 inst_Module70();
    Module40 inst_Module40();
    Module29 inst_Module29();
endmodule
