module rootModule_1_1_0();
    rootModule_1_1_0_0 inst_0();
    rootModule_1_1_0_1 inst_1();
endmodule
