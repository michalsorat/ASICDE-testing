module Module80();
    Module89 inst_Module89();
    Module82 inst_Module82();
    Module97 inst_Module97();
    Module92 inst_Module92();
    Module88 inst_Module88();
endmodule
