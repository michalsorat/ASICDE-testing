module Module45();
    Module59 inst_Module59();
    Module46 inst_Module46();
endmodule
