module rootModule_sb0_0_sb1_1_sb2_0_sb3_2_sb4_1();
endmodule
