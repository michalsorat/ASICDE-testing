module rootModule_2_0_0_0();
    rootModule_2_0_0_0_0 inst_0();
    rootModule_2_0_0_0_1 inst_1();
endmodule
