module Module12();
    Module94 inst_Module94();
endmodule
