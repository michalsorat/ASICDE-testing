module rootModule_sub_0_0_sub_1_2();
    rootModule_sub_0_0_sub_1_2_sub_2_0 inst_0();
    rootModule_sub_0_0_sub_1_2_sub_2_1 inst_1();
endmodule
