module rootModule_sub_0_0();
    rootModule_sub_0_0_sub_1_0 inst_0();
endmodule
