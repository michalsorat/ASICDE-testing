module rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_0 inst_0();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_1 inst_1();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_2 inst_2();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_3 inst_3();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_4 inst_4();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_5 inst_5();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_6 inst_6();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_7 inst_7();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_8 inst_8();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_2_sw18_7_sw19_9 inst_9();
endmodule
