module rootModule_2_2_1();
    rootModule_2_2_1_0 inst_0();
endmodule
