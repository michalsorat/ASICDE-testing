module rootModule_1_0_0_0_1();
endmodule
