module rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0();
    rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0 inst_0();
endmodule
