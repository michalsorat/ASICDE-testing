module rootModule_1_0_2_0();
    rootModule_1_0_2_0_0 inst_0();
endmodule
