module Module90();
    Module94 inst_Module94();
    Module92 inst_Module92();
endmodule
