module Module33();
    Module94 inst_Module94();
    Module61 inst_Module61();
    Module69 inst_Module69();
endmodule
