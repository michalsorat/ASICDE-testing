module Module70();
    Module88 inst_Module88();
    Module81 inst_Module81();
    Module78 inst_Module78();
    Module93 inst_Module93();
endmodule
