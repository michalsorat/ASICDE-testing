module rootModule_1_1_1_1();
    rootModule_1_1_1_1_0 inst_0();
endmodule
