module rootModule1000();
    rootModule1000_sf0_0 inst_0();
endmodule
