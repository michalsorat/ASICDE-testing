module Module86();
    Module95 inst_Module95();
    Module98 inst_Module98();
endmodule
