module rootModule_sub_0_0_sub_1_0_sub_2_2();
    rootModule_sub_0_0_sub_1_0_sub_2_2_sub_3_0 inst_0();
    rootModule_sub_0_0_sub_1_0_sub_2_2_sub_3_1 inst_1();
endmodule
