module rootModule1000_se0_0_se1_0();
    rootModule1000_se0_0_se1_0_se2_0 inst_0();
endmodule
