module rootModule_1_1_1_1_0();
endmodule
