module Module25();
    Module27 inst_Module27();
    Module30 inst_Module30();
    Module51 inst_Module51();
    Module82 inst_Module82();
    Module63 inst_Module63();
endmodule
