module Module41();
    Module93 inst_Module93();
    Module52 inst_Module52();
    Module70 inst_Module70();
    Module63 inst_Module63();
    Module43 inst_Module43();
endmodule
