module rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_1_sf7_3_sf8_0();
    rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_1_sf7_3_sf8_0_sf9_0 inst_0();
    rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_1_sf7_3_sf8_0_sf9_1 inst_1();
    rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_1_sf7_3_sf8_0_sf9_2 inst_2();
    rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_1_sf7_3_sf8_0_sf9_3 inst_3();
    rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_1_sf7_3_sf8_0_sf9_4 inst_4();
endmodule
