module rootModule();
    rootModule_sb0_0 inst_0();
    rootModule_sb0_1 inst_1();
    rootModule_sb0_2 inst_2();
endmodule
