module rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_0 inst_0();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_1 inst_1();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_2 inst_2();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_3 inst_3();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_4 inst_4();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_5 inst_5();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_6 inst_6();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_7 inst_7();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_8 inst_8();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_9 inst_9();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_10 inst_10();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_11 inst_11();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_12 inst_12();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_13 inst_13();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_1_s28_13_s29_14 inst_14();
endmodule
