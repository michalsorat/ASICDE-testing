module rootModule_sb0_0_sb1_0_sb2_1_sb3_2_sb4_0();
endmodule
