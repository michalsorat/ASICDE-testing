module rootModule_1_1_1_2_1();
endmodule
