module Module21();
    Module25 inst_Module25();
    Module48 inst_Module48();
    Module80 inst_Module80();
    Module69 inst_Module69();
endmodule
