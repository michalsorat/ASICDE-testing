module rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0 inst_0();
endmodule
