module rootModule1000();
    rootModule1000_s0_0 inst_0();
endmodule
