module rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_1_sc9_2();
endmodule
