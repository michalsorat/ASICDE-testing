module rootModule_1_1_0_1_0();
endmodule
