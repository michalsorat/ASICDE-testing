module rootModule_0_0();
    rootModule_0_0_0 inst_0();
endmodule
