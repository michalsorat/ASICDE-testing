module rootModule_sub0_0_sub1_1_sub2_2_sub3_2_sub4_0();
endmodule
