module Module23();
    Module47 inst_Module47();
    Module82 inst_Module82();
    Module89 inst_Module89();
    Module48 inst_Module48();
    Module66 inst_Module66();
endmodule
