module rootModule_sub0_0_sub1_0_sub2_0_sub3_1_sub4_2();
    rootModule_sub0_0_sub1_0_sub2_0_sub3_1_sub4_2_sub5_0 inst_0();
    rootModule_sub0_0_sub1_0_sub2_0_sub3_1_sub4_2_sub5_1 inst_1();
    rootModule_sub0_0_sub1_0_sub2_0_sub3_1_sub4_2_sub5_2 inst_2();
endmodule
