module rootModule_sub0_0_sub1_1_sub2_1_sub3_2();
    rootModule_sub0_0_sub1_1_sub2_1_sub3_2_sub4_0 inst_0();
    rootModule_sub0_0_sub1_1_sub2_1_sub3_2_sub4_1 inst_1();
    rootModule_sub0_0_sub1_1_sub2_1_sub3_2_sub4_2 inst_2();
endmodule
