module Module22();
    Module28 inst_Module28();
    Module56 inst_Module56();
endmodule
