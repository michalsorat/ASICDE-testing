module rootModule_1_1_2_2_1();
endmodule
