module Module10();
    Module41 inst_Module41();
    Module14 inst_Module14();
    Module68 inst_Module68();
    Module43 inst_Module43();
    Module17 inst_Module17();
endmodule
