module rootModule1000_s0_0_s1_0_s2_0();
    rootModule1000_s0_0_s1_0_s2_0_s3_0 inst_0();
endmodule
