module Module87();
    Module92 inst_Module92();
endmodule
