module Module9();
    Module93 inst_Module93();
    Module96 inst_Module96();
endmodule
