module Module7();
    Module74 inst_Module74();
    Module48 inst_Module48();
endmodule
