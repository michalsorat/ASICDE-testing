module Module68();
    Module92 inst_Module92();
    Module83 inst_Module83();
    Module84 inst_Module84();
    Module76 inst_Module76();
endmodule
