module Module88();
    Module99 inst_Module99();
    Module96 inst_Module96();
    Module98 inst_Module98();
endmodule
