module rootModule();
    rootModule_sub_0_0 inst_0();
endmodule
