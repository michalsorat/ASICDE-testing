module rootModule_0_0_0_1_1();
endmodule
