module rootModule();
    rootModule_sub_0_0 inst_0();
    rootModule_sub_0_1 inst_1();
endmodule
