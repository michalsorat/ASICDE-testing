module rootModule_sb0_0_sb1_2_sb2_2_sb3_1();
    rootModule_sb0_0_sb1_2_sb2_2_sb3_1_sb4_0 inst_0();
    rootModule_sb0_0_sb1_2_sb2_2_sb3_1_sb4_1 inst_1();
    rootModule_sb0_0_sb1_2_sb2_2_sb3_1_sb4_2 inst_2();
endmodule
