module rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0();
    rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0 inst_0();
endmodule
