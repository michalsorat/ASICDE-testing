module Module89();
    Module96 inst_Module96();
    Module90 inst_Module90();
    Module97 inst_Module97();
    Module93 inst_Module93();
endmodule
