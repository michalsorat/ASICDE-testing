module rootModule300_sw0_0_sw1_0();
    rootModule300_sw0_0_sw1_0_sw2_0 inst_0();
endmodule
