module rootModule_2_0_0_0_1();
endmodule
