module rootModule_sb0_1_sb1_0_sb2_2_sb3_1_sb4_0();
endmodule
