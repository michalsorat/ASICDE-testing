module rootModule_2_1_1_1_2();
endmodule
