module rootModule();
    rootModule_sb0_0 inst_0();
endmodule
