module rootModule();
    rootModule_sub0_0 inst_0();
endmodule
