module rootModule_1_1_2_0_0();
endmodule
