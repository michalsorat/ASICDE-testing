module Module95();
    Module99 inst_Module99();
endmodule
