module rootModule_sb0_2_sb1_0_sb2_1_sb3_1_sb4_2();
endmodule
