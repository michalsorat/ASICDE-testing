module rootModule_2_2_2_0_0();
endmodule
