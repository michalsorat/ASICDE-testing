module rootModule_2_0_1_1_1();
endmodule
