module rootModule_sg0_0_sg1_0_sg2_0_sg3_0_sg4_0_sg5_0_sg6_0_sg7_1_sg8_3_sg9_1();
endmodule
