module rootModule_1_0_2_0_0();
endmodule
