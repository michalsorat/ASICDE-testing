module Module20();
    Module96 inst_Module96();
    Module82 inst_Module82();
endmodule
