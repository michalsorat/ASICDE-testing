module rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_1();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_1_sd8_0 inst_0();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_1_sd8_1 inst_1();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_1_sd8_2 inst_2();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_1_sd8_3 inst_3();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_1_sd8_4 inst_4();
endmodule
