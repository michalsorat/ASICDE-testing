module rootModule_2_2();
    rootModule_2_2_0 inst_0();
    rootModule_2_2_1 inst_1();
    rootModule_2_2_2 inst_2();
endmodule
