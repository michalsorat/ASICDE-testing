module rootModule1000();
    rootModule1000_sc0_0 inst_0();
endmodule
