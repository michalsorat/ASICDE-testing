module Module6();
    Module33 inst_Module33();
endmodule
