module rootModule_0_0_0_1_2();
endmodule
