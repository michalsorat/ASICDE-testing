module Module78();
    Module96 inst_Module96();
endmodule
