module Module50();
    Module76 inst_Module76();
    Module85 inst_Module85();
    Module95 inst_Module95();
    Module79 inst_Module79();
    Module96 inst_Module96();
endmodule
