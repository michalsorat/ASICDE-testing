module rootModule1000_s0_0_s1_0_s2_0_s3_0_s4_0_s5_0_s6_0_s7_0_s8_0_s9_0_s10_0_s11_0_s12_0_s13_0_s14_0_s15_0_s16_0_s17_0_s18_0_s19_0_s20_0_s21_0_s22_0_s23_0_s24_0_s25_0_s26_0_s27_3_s28_14_s29_11();
endmodule
