module rootModule_1_0_1_0();
    rootModule_1_0_1_0_0 inst_0();
endmodule
