module rootModule1000_sd0_0();
    rootModule1000_sd0_0_sd1_0 inst_0();
endmodule
