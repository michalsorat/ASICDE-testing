module rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_1_sb18_3_sb19_4();
endmodule
