module Module65();
    Module84 inst_Module84();
    Module95 inst_Module95();
    Module86 inst_Module86();
endmodule
