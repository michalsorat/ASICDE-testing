module rootModule_sb0_1_sb1_1_sb2_0_sb3_0();
    rootModule_sb0_1_sb1_1_sb2_0_sb3_0_sb4_0 inst_0();
    rootModule_sb0_1_sb1_1_sb2_0_sb3_0_sb4_1 inst_1();
    rootModule_sb0_1_sb1_1_sb2_0_sb3_0_sb4_2 inst_2();
endmodule
