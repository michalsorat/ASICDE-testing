module Module71();
    Module85 inst_Module85();
    Module73 inst_Module73();
    Module92 inst_Module92();
endmodule
