module rootModule();
    rootModule_sw0_0 inst_0();
endmodule
