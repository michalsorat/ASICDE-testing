module Module36();
    Module38 inst_Module38();
    Module79 inst_Module79();
endmodule
