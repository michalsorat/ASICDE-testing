module rootModule();
    rootModule_sg0_0 inst_0();
endmodule
