module Module77();
    Module90 inst_Module90();
    Module81 inst_Module81();
    Module84 inst_Module84();
    Module93 inst_Module93();
endmodule
