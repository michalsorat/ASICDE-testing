module Module2();
    Module69 inst_Module69();
endmodule
