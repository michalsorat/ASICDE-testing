module rootModule_0_0_0_1_0();
endmodule
