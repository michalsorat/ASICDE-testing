module Module48();
    Module71 inst_Module71();
    Module51 inst_Module51();
endmodule
