module rootModule_sb0_2();
    rootModule_sb0_2_sb1_0 inst_0();
    rootModule_sb0_2_sb1_1 inst_1();
endmodule
