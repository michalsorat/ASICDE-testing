module Module74();
    Module78 inst_Module78();
    Module81 inst_Module81();
    Module82 inst_Module82();
    Module95 inst_Module95();
    Module92 inst_Module92();
endmodule
