module rootModule_1_0_2_1_0();
endmodule
