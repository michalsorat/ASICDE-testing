module rootModule_sub0_0_sub1_0_sub2_1_sub3_0_sub4_0();
endmodule
