module rootModule_2_0_1_1_2();
endmodule
