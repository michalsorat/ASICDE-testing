module Module97();
    Module99 inst_Module99();
endmodule
