module rootModule_sb0_1_sb1_2_sb2_1_sb3_2_sb4_0();
endmodule
