module Module76();
    Module97 inst_Module97();
    Module93 inst_Module93();
    Module85 inst_Module85();
endmodule
