module rootModule_sb0_1_sb1_1_sb2_0_sb3_1_sb4_0();
endmodule
