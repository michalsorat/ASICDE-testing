module rootModule_1_1_1_2_0();
endmodule
