module rootModule_0_0_0_1();
    rootModule_0_0_0_1_0 inst_0();
    rootModule_0_0_0_1_1 inst_1();
    rootModule_0_0_0_1_2 inst_2();
endmodule
