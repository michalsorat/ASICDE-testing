module rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_1_se7_1_se8_2_se9_1();
endmodule
