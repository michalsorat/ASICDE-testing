module rootModule_sub_0_1();
    rootModule_sub_0_1_sub_1_0 inst_0();
    rootModule_sub_0_1_sub_1_1 inst_1();
endmodule
