module Module31();
    Module63 inst_Module63();
    Module34 inst_Module34();
    Module42 inst_Module42();
    Module68 inst_Module68();
    Module47 inst_Module47();
endmodule
