module Module82();
    Module95 inst_Module95();
    Module97 inst_Module97();
    Module88 inst_Module88();
    Module96 inst_Module96();
    Module98 inst_Module98();
endmodule
