module Module64();
    Module95 inst_Module95();
    Module73 inst_Module73();
endmodule
