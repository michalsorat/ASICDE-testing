module rootModule_sb0_1_sb1_0_sb2_1_sb3_0_sb4_0();
endmodule
