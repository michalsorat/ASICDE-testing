module Module18();
    Module23 inst_Module23();
    Module60 inst_Module60();
    Module68 inst_Module68();
endmodule
