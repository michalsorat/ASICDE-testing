module rootModule1000_sc0_0();
    rootModule1000_sc0_0_sc1_0 inst_0();
endmodule
