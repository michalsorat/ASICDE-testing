module Module13();
    Module43 inst_Module43();
    Module28 inst_Module28();
endmodule
