module rootModule_sub0_0_sub1_2_sub2_0_sub3_1_sub4_2();
endmodule
