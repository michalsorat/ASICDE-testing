module Module67();
    Module71 inst_Module71();
    Module76 inst_Module76();
    Module80 inst_Module80();
endmodule
