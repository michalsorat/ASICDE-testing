module rootModule_sb0_0_sb1_0_sb2_1();
    rootModule_sb0_0_sb1_0_sb2_1_sb3_0 inst_0();
    rootModule_sb0_0_sb1_0_sb2_1_sb3_1 inst_1();
    rootModule_sb0_0_sb1_0_sb2_1_sb3_2 inst_2();
endmodule
