module rootModule_sub0_0_sub1_0_sub2_2_sub3_1();
    rootModule_sub0_0_sub1_0_sub2_2_sub3_1_sub4_0 inst_0();
endmodule
