module rootModule_2_1_1_2_0();
endmodule
