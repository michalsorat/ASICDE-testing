module rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_3_sw8_1();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_3_sw8_1_sw9_0 inst_0();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_3_sw8_1_sw9_1 inst_1();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_3_sw8_1_sw9_2 inst_2();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_3_sw8_1_sw9_3 inst_3();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_3_sw8_1_sw9_4 inst_4();
endmodule
