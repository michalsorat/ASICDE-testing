module Module40();
    Module82 inst_Module82();
    Module52 inst_Module52();
    Module99 inst_Module99();
    Module44 inst_Module44();
    Module91 inst_Module91();
endmodule
