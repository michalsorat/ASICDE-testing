module rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0_sw7_0_sw8_0_sw9_0_sw10_0_sw11_0_sw12_0_sw13_0_sw14_0_sw15_0_sw16_0_sw17_1_sw18_4_sw19_3();
endmodule
