module rootModule1000_sf0_0();
    rootModule1000_sf0_0_sf1_0 inst_0();
endmodule
