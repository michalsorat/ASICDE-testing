module rootModule_2_2_2();
    rootModule_2_2_2_0 inst_0();
endmodule
