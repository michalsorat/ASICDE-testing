module Module29();
    Module98 inst_Module98();
endmodule
