module Module19();
    Module39 inst_Module39();
    Module56 inst_Module56();
endmodule
