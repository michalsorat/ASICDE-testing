module rootModule_sub0_0_sub1_1_sub2_2_sub3_1_sub4_2();
endmodule
