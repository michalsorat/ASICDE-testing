module rootModule_sub0_0_sub1_1_sub2_2_sub3_0_sub4_1();
endmodule
