module Module66();
    Module70 inst_Module70();
    Module71 inst_Module71();
endmodule
