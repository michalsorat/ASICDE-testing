module Module75();
    Module85 inst_Module85();
    Module84 inst_Module84();
endmodule
