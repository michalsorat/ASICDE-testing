module rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_2();
    rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_2_sc9_0 inst_0();
    rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_2_sc9_1 inst_1();
    rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_2_sc9_2 inst_2();
    rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_2_sc9_3 inst_3();
    rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0_sc6_1_sc7_0_sc8_2_sc9_4 inst_4();
endmodule
