module rootModule_sb0_2_sb1_0_sb2_1_sb3_2();
    rootModule_sb0_2_sb1_0_sb2_1_sb3_2_sb4_0 inst_0();
    rootModule_sb0_2_sb1_0_sb2_1_sb3_2_sb4_1 inst_1();
    rootModule_sb0_2_sb1_0_sb2_1_sb3_2_sb4_2 inst_2();
endmodule
