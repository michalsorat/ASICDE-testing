module Module73();
    Module96 inst_Module96();
    Module99 inst_Module99();
endmodule
