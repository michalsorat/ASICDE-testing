module rootModule_sub_0_1_sub_1_1_sub_2_0_sub_3_0_sub_4_2();
endmodule
