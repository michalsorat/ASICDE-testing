module rootModule_2_0_1();
    rootModule_2_0_1_0 inst_0();
    rootModule_2_0_1_1 inst_1();
endmodule
