module rootModule_sub_0_0_sub_1_0_sub_2_2_sub_3_1_sub_4_0();
endmodule
