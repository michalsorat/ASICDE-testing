module Module60();
    Module61 inst_Module61();
    Module76 inst_Module76();
    Module97 inst_Module97();
endmodule
