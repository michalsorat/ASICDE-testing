module rootModule_0();
    rootModule_0_0 inst_0();
endmodule
