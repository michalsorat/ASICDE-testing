module rootModule_sub_0_1_sub_1_1();
    rootModule_sub_0_1_sub_1_1_sub_2_0 inst_0();
endmodule
