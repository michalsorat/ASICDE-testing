module Module11();
    Module36 inst_Module36();
    Module83 inst_Module83();
endmodule
