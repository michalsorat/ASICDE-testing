module rootModule_1();
    rootModule_1_0 inst_0();
    rootModule_1_1 inst_1();
endmodule
