module Module83();
    Module91 inst_Module91();
    Module92 inst_Module92();
endmodule
