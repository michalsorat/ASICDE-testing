module Module27();
    Module42 inst_Module42();
    Module51 inst_Module51();
    Module36 inst_Module36();
    Module67 inst_Module67();
    Module85 inst_Module85();
endmodule
