module rootModule_2_2_1_0();
    rootModule_2_2_1_0_0 inst_0();
    rootModule_2_2_1_0_1 inst_1();
    rootModule_2_2_1_0_2 inst_2();
endmodule
