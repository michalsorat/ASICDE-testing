module Module28();
    Module81 inst_Module81();
    Module94 inst_Module94();
    Module96 inst_Module96();
    Module83 inst_Module83();
    Module64 inst_Module64();
endmodule
