module rootModule_2_1_1();
    rootModule_2_1_1_0 inst_0();
    rootModule_2_1_1_1 inst_1();
    rootModule_2_1_1_2 inst_2();
endmodule
