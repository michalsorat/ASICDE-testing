module rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0();
    rootModule1000_sc0_0_sc1_0_sc2_0_sc3_0_sc4_0_sc5_0 inst_0();
endmodule
