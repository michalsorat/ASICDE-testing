module rootModule_2_0_1_0_2();
endmodule
