module Module49();
    Module79 inst_Module79();
    Module68 inst_Module68();
    Module93 inst_Module93();
    Module87 inst_Module87();
    Module76 inst_Module76();
endmodule
