module Module17();
    Module31 inst_Module31();
endmodule
