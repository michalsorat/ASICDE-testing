module rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0 inst_0();
    rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_1 inst_1();
endmodule
