module rootModule1000_sf0_0_sf1_0_sf2_0_sf3_0_sf4_0_sf5_0_sf6_2_sf7_1_sf8_2_sf9_3();
endmodule
