module rootModule1000_sd0_0_sd1_0_sd2_0_sd3_0_sd4_0_sd5_0_sd6_0_sd7_4_sd8_4_sd9_0();
endmodule
