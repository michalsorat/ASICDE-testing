module Module37();
    Module92 inst_Module92();
    Module91 inst_Module91();
endmodule
