module rootModule1000_se0_0_se1_0_se2_0_se3_0_se4_0_se5_0_se6_0_se7_2_se8_1_se9_3();
endmodule
