module rootModule_sb0_0_sb1_0_sb2_0();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0 inst_0();
endmodule
