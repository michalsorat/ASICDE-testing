module rootModule_1_0_2_1_1();
endmodule
