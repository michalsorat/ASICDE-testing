module rootModule_sub0_0();
    rootModule_sub0_0_sub1_0 inst_0();
    rootModule_sub0_0_sub1_1 inst_1();
    rootModule_sub0_0_sub1_2 inst_2();
endmodule
