module Module91();
    Module97 inst_Module97();
endmodule
