module rootModule_sw0_0_sw1_0();
    rootModule_sw0_0_sw1_0_sw2_0 inst_0();
endmodule
