module rootModule_sb0_0_sb1_0_sb2_1_sb3_1_sb4_1();
endmodule
