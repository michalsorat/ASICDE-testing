module rootModule_sub0_0_sub1_1_sub2_0_sub3_0_sub4_0();
endmodule
