module rootModule_sub0_0_sub1_2_sub2_1();
    rootModule_sub0_0_sub1_2_sub2_1_sub3_0 inst_0();
endmodule
