module Module43();
    Module55 inst_Module55();
    Module86 inst_Module86();
endmodule
