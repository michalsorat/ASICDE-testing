module rootModule_1_0_2_1_2();
endmodule
