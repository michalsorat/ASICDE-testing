module Module98();
    Module99 inst_Module99();
endmodule
