module Module69();
    Module74 inst_Module74();
    Module80 inst_Module80();
    Module79 inst_Module79();
    Module96 inst_Module96();
    Module83 inst_Module83();
endmodule
