module rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_1_sw7_1_sw8_2_sw9_0();
endmodule
