module rootModule300();
    rootModule300_sw0_0 inst_0();
endmodule
