module Module0();
    Module7 inst_Module7();
    Module1 inst_Module1();
    Module84 inst_Module84();
    Module83 inst_Module83();
endmodule
