module Module4();
    Module69 inst_Module69();
    Module32 inst_Module32();
    Module38 inst_Module38();
endmodule
