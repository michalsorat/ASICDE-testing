module Module94();
    Module95 inst_Module95();
    Module96 inst_Module96();
    Module98 inst_Module98();
    Module99 inst_Module99();
    Module97 inst_Module97();
endmodule
