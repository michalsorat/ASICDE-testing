module Module92();
    Module99 inst_Module99();
    Module97 inst_Module97();
endmodule
