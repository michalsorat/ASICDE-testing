module Module63();
    Module97 inst_Module97();
endmodule
