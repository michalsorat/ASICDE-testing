module Module42();
    Module62 inst_Module62();
    Module92 inst_Module92();
endmodule
