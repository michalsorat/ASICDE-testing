module Module8();
    Module80 inst_Module80();
endmodule
