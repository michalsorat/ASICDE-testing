module Module39();
    Module86 inst_Module86();
    Module60 inst_Module60();
    Module46 inst_Module46();
endmodule
