module Module35();
    Module41 inst_Module41();
    Module95 inst_Module95();
    Module92 inst_Module92();
    Module66 inst_Module66();
    Module39 inst_Module39();
endmodule
