module rootModule_0_0_0_0_0();
endmodule
