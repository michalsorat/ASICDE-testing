module Module79();
    Module99 inst_Module99();
endmodule
