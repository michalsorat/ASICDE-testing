module rootModule1000();
    rootModule1000_se0_0 inst_0();
endmodule
