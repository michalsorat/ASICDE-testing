module rootModule_1_1_2_0();
    rootModule_1_1_2_0_0 inst_0();
endmodule
