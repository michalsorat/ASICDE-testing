module Module14();
    Module35 inst_Module35();
endmodule
