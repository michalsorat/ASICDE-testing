module rootModule1000();
    rootModule1000_sd0_0 inst_0();
endmodule
