module rootModule_2_1_1_0_0();
endmodule
