module Module44();
    Module74 inst_Module74();
    Module46 inst_Module46();
    Module53 inst_Module53();
    Module89 inst_Module89();
    Module64 inst_Module64();
endmodule
