module rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0 inst_0();
    rootModule300_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_1 inst_1();
endmodule
