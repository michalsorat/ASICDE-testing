module Module99();
endmodule
