module rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0();
    rootModule_sw0_0_sw1_0_sw2_0_sw3_0_sw4_0_sw5_0_sw6_0 inst_0();
endmodule
