module Module53();
    Module96 inst_Module96();
endmodule
