module rootModule_0_0_0_0_1();
endmodule
