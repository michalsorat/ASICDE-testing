module Module47();
    Module59 inst_Module59();
    Module73 inst_Module73();
endmodule
