module rootModule_1_0_1_0_0();
endmodule
