module Module84();
    Module97 inst_Module97();
    Module96 inst_Module96();
    Module99 inst_Module99();
    Module94 inst_Module94();
endmodule
