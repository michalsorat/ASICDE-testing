module rootModule();
    Module73 inst_Module73();
    Module18 inst_Module18();
    Module65 inst_Module65();
    Module10 inst_Module10();
    Module12 inst_Module12();
endmodule
