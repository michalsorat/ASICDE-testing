module rootModule_2_1_1_1_1();
endmodule
