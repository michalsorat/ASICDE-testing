module rootModule_sb0_1();
    rootModule_sb0_1_sb1_0 inst_0();
    rootModule_sb0_1_sb1_1 inst_1();
    rootModule_sb0_1_sb1_2 inst_2();
endmodule
