module rootModule_sub0_0_sub1_0_sub2_0_sub3_2();
    rootModule_sub0_0_sub1_0_sub2_0_sub3_2_sub4_0 inst_0();
    rootModule_sub0_0_sub1_0_sub2_0_sub3_2_sub4_1 inst_1();
    rootModule_sub0_0_sub1_0_sub2_0_sub3_2_sub4_2 inst_2();
endmodule
