module Module59();
    Module91 inst_Module91();
    Module89 inst_Module89();
    Module87 inst_Module87();
endmodule
