module Module85();
    Module89 inst_Module89();
endmodule
