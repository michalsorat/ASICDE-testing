module Module46();
    Module70 inst_Module70();
    Module69 inst_Module69();
    Module87 inst_Module87();
endmodule
