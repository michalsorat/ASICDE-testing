module Module54();
    Module92 inst_Module92();
    Module97 inst_Module97();
    Module61 inst_Module61();
    Module86 inst_Module86();
    Module95 inst_Module95();
endmodule
