module rootModule();
    rootModule_0 inst_0();
    rootModule_1 inst_1();
    rootModule_2 inst_2();
endmodule
