module Module15();
    Module90 inst_Module90();
    Module69 inst_Module69();
    Module65 inst_Module65();
    Module34 inst_Module34();
endmodule
