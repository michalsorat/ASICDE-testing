module Module5();
    Module87 inst_Module87();
    Module18 inst_Module18();
    Module53 inst_Module53();
    Module54 inst_Module54();
    Module27 inst_Module27();
endmodule
