module Module72();
    Module93 inst_Module93();
endmodule
