module rootModule_sub0_0_sub1_0_sub2_2_sub3_2_sub4_2();
endmodule
