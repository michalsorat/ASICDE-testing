module rootModule_1_1_2_1_1();
endmodule
