module rootModule_2_1_0();
    rootModule_2_1_0_0 inst_0();
endmodule
