module rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_0 inst_0();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_1 inst_1();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_2 inst_2();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_3 inst_3();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_4 inst_4();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_5 inst_5();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_6 inst_6();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_7 inst_7();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_8 inst_8();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0_sb7_0_sb8_0_sb9_0_sb10_0_sb11_0_sb12_0_sb13_0_sb14_0_sb15_0_sb16_0_sb17_0_sb18_4_sb19_9 inst_9();
endmodule
