module rootModule1000_s0_0_s1_0();
    rootModule1000_s0_0_s1_0_s2_0 inst_0();
endmodule
