module Module55();
    Module57 inst_Module57();
    Module84 inst_Module84();
endmodule
