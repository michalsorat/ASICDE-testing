module rootModule_2_2_2_0_1();
endmodule
