module rootModule_sub_0_0_sub_1_1_sub_2_2_sub_3_1_sub_4_2();
    rootModule_sub_0_0_sub_1_1_sub_2_2_sub_3_1_sub_4_2_sub_5_0 inst_0();
    rootModule_sub_0_0_sub_1_1_sub_2_2_sub_3_1_sub_4_2_sub_5_1 inst_1();
    rootModule_sub_0_0_sub_1_1_sub_2_2_sub_3_1_sub_4_2_sub_5_2 inst_2();
endmodule
