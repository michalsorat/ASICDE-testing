module rootModule_1_1_1_2();
    rootModule_1_1_1_2_0 inst_0();
    rootModule_1_1_1_2_1 inst_1();
endmodule
