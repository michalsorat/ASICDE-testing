module rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0();
    rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0_sb5_0_sb6_0 inst_0();
endmodule
