module Module61();
    Module97 inst_Module97();
endmodule
