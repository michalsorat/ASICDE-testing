module rootModule_sb0_2_sb1_1_sb2_1();
endmodule
