module Module96();
    Module99 inst_Module99();
endmodule
