module Module62();
    Module76 inst_Module76();
endmodule
