module Module52();
    Module97 inst_Module97();
    Module54 inst_Module54();
    Module63 inst_Module63();
    Module85 inst_Module85();
    Module82 inst_Module82();
endmodule
