module rootModule_sb0_0_sb1_0_sb2_0_sb3_0_sb4_0();
endmodule
