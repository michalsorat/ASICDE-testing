module rootModule_2_1_1_2_1();
endmodule
